
`ifndef JTAG_AGENT_SV
`define JTAG_AGENT_SV

class jtag_agent extends uvm_agent;
    `uvm_component_utils(jtag_agent)
    
    jtag_driver driver;
    jtag_monitor monitor;
    jtag_sequencer sequencer;
    jtag_config cfg;
    
    function new(string name, uvm_component parent);
        super.new(name, parent);
    endfunction
    
    function void build_phase(uvm_phase phase);
        super.build_phase(phase);
        
        if(!uvm_config_db#(jtag_config)::get(this, "", "cfg", cfg)) begin
            `uvm_fatal("NOCFG", "Config object not set")
        end
        
        monitor = jtag_monitor::type_id::create("monitor", this);
        
        if(cfg.active_passive == UVM_ACTIVE) begin
            driver = jtag_driver::type_id::create("driver", this);
            sequencer = jtag_sequencer::type_id::create("sequencer", this);
        end
    endfunction
    
    function void connect_phase(uvm_phase phase);
        super.connect_phase(phase);
        
        if(cfg.active_passive == UVM_ACTIVE) begin
            driver.seq_item_port.connect(sequencer.seq_item_export);
        end
        
        // Connect virtual interface to driver and monitor
        uvm_config_db#(virtual jtag_if)::set(this, "driver", "vif", cfg.vif);
        uvm_config_db#(virtual jtag_if)::set(this, "monitor", "vif", cfg.vif);
        uvm_config_db#(jtag_config)::set(this, "driver", "cfg", cfg);
        uvm_config_db#(jtag_config)::set(this, "monitor", "cfg", cfg);
    endfunction
endclass

`endif //JTAG_AGENT_SV
